module bttn (
    input [3:0] bttns,
    output [3:0] pmod
);

assign bttns = pmod;

endmodule

module ledTest2 (
    input
)
// Buton verisi eklenecek TO-DO
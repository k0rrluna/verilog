module andSixTGateTB();
    reg [15:0] A_i;
    reg [15:0] B_i;
    wire [15:0] Y_o;

    andSixTGate uut(
        .A_i(A_i),
        .B_i(B_i),
        .Y_o(Y_o)
);

initial begin
    $dumpfile("andSixTGate.vcd");
    $dumpvars;
    A_i = 16'b0000_0000_0000_0000; B_i = 16'b0000_0000_0000_0000; #10;
    A_i = 16'b0000_0000_0000_0000; B_i = 16'b0000_0000_0000_0001; #10;
    A_i = 16'b0000_0000_0000_0001; B_i = 16'b0000_0000_0000_0001; #10;
    A_i = 16'b0000_0000_0100_0000; B_i = 16'b0000_0000_0000_0000; #10;
    A_i = 16'b0000_0000_0100_0000; B_i = 16'b0000_0000_0100_0000; #10;
    A_i = 16'b0000_0000_0000_0000; B_i = 16'b0000_0010_0000_0000; #10;
    A_i = 16'b0000_0010_0000_0000; B_i = 16'b0000_0010_0000_0000; #10;
    A_i = 16'b1111_1111_1111_1111; B_i = 16'b1111_1111_1111_1111; #10;
    $finish;
end

endmodule
